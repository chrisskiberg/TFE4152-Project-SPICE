* Check OP

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../models/ptm_130.spi
.include ../../lib/SUN_TR_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-20 reltol=1e-8 abstol=1e-10

*----------------------------------------------------------------
* PARAMETERS - must change for correct operating region
*----------------------------------------------------------------
.param VDD_param = 1.5

.param BIAS1 = 0.72
.param BIAS2 = 0.44
.param VSTORE_param = 1.0

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------

V1 VDD 0 dc VDD_param
V2 VSS 0 dc 0

VBIAS1 VBIAS1 0 dc BIAS1
VBIAS2 VBIAS2 0 dc BIAS2	

VSTORE VSTORE 0 dc VSTORE_param

*----------------------------------------------------------------
* RAMP
*----------------------------------------------------------------
VRAMP VRAMP 0 dc 1.3

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include comparator_test.cir

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------

X1 VSTORE VRAMP VBIAS1 VBIAS2 VDD VSS VCMP_OUT COMP

*----------------------------------------------------------------
* Analysis 
*----------------------------------------------------------------
.op

