.SUBCKT PIXEL_SENSOR VBIAS1 VBIAS2 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR
XC1 VSTORE VRAMP VBIAS1 VBIAS2 VDD VSS VCMP_OUT COMP
XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS


.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS
XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL
.ENDS


.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS

.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

* Capacitor to model gate-source capacitance
C1 VSTORE VSS 100f
Rleak VSTORE VSS 100T

* Switch to reset voltage on capacitor
BR1 VRESET VSTORE I=V(ERASE)*V(VRESET,VSTORE)/1k

* Switch to expose pixel
BR2 VPG VSTORE I=V(EXPOSE)*V(VSTORE,VPG)/1k

* Model photocurrent
Rphoto VPG VSS 1G
.ENDS

.SUBCKT COMP VSTORE VRAMP VBIAS1 VBIAS2 VDD VSS VCMP_OUT
MCML VCMOL VCMOL VDD VDD pmos L=0.5u W=0.5u 
MCMR VCMOR VCMOL VDD VDD pmos L=0.5u W=0.5u

MDPR VCMOR VRAMP VDPCI VSS nmos L=0.15u W=0.65u
MDPL VCMOL VSTORE VDPCI VSS nmos L=0.15u W=0.65u 

MDPC VDPCI VBIAS1 VSS VSS nmos L=0.8u W=0.13u 

MIP1 VIP1 VCMOR VDD VDD pmos W=0.65u L=0.13u
MIN1 VIP1 VBIAS2 VSS VSS nmos W=0.65u L=0.13u

MIP2 VCMP_OUT VIP1 VDD VDD pmos W=0.65u L=0.13u
MIN2 VCMP_OUT VIP1 VSS VSS nmos W=0.65u L=0.13u
.ENDS