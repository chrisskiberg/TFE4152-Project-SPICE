.subckt COMP VSTORE VRAMP VBIAS1 VBIAS2 VDD VSS VCMP_OUT
MCML VCMOL VCMOL VDD VDD pmos L=0.5u W=0.5u 
MCMR VCMOR VCMOL VDD VDD pmos L=0.5u W=0.5u

MDPR VCMOR VRAMP VDPCI VSS nmos L=0.15u W=0.65u
MDPL VCMOL VSTORE VDPCI VSS nmos L=0.15u W=0.65u 

MDPC VDPCI VBIAS1 VSS VSS nmos L=0.8u W=0.13u 

MIP1 VIP1 VCMOR VDD VDD pmos W=0.65u L=0.13u
MIN1 VIP1 VBIAS2 VSS VSS nmos W=0.65u L=0.13u

MIP2 VCMP_OUT VIP1 VDD VDD pmos W=0.65u L=0.13u
MIN2 VCMP_OUT VIP1 VSS VSS nmos W=0.65u L=0.13u
.ends